/*************************************************************************
*
* Copyright © Microsoft Corporation. All rights reserved.
* Copyright © Broadcom Inc. All rights reserved.
* Licensed under the MIT License.
*
*************************************************************************/
module CR_TIE_CELL(ob, o);
   output wire ob ;
   output wire o;


   assign      o  = 1'b1;
   assign      ob = 1'b0;
   
endmodule 

/*************************************************************************
*
* Copyright � Microsoft Corporation. All rights reserved.
* Copyright � Broadcom Inc. All rights reserved.
* Licensed under the MIT License.
*
*************************************************************************/









`ifndef __CR_HUF_COMP_VH
`define __CR_HUF_COMP_VH


`include "cr_huf_comp_regs.vh"
`include "cr_huf_comp_regsPKG.svp"
`include "cr_huf_comp_regfilePKG.svp"


`define MAX(a,b) \
    (((a)>(b))?(a):(b))
`define MIN(a,b) \
    (((a)<(b))?(a):(b))
`define LOG_VEC(a) `MAX(0, ($clog2(a)-1)):0
`define ROUND_UP_DIV(a,b) \
    ((a%b)==0 ? (a/b) : (a/b)+1)


`define CLK_GATE   



`define CREOLE_HC_SHORT_DAT_WIDTH `N_SHRT_SYM_WIDTH
`define CREOLE_HC_SHORT_CNT_WIDTH 3
`define CREOLE_HC_SHORT_FREQ_WIDTH 16
`define CREOLE_HC_LONG_DAT_WIDTH `N_LONG_SYM_WIDTH
`define CREOLE_HC_LONG_CNT_WIDTH 1
`define CREOLE_HC_LONG_FREQ_WIDTH 14
`define CREOLE_HC_SHORT_NUM_MAX_SYM_USED 576
`define CREOLE_HC_SHORT_SYM_ADDR_WIDTH $clog2(`CREOLE_HC_SHORT_NUM_MAX_SYM_USED)
`define CREOLE_HC_LONG_NUM_MAX_SYM_USED 248
`define CREOLE_HC_LONG_SYM_ADDR_WIDTH $clog2(`CREOLE_HC_LONG_NUM_MAX_SYM_USED)
`define CREOLE_HC_SEQID_NUM 10
`define CREOLE_HC_SEQID_WIDTH 4
`define CREOLE_HC_SYMBOL_QUEUE_WIDTH 75 
`define CREOLE_HC_PHT_WIDTH 60
`define CREOLE_HC_PHT_ADDR_WIDTH 6
`define CREOLE_HC_HDR_WIDTH 64
`define CREOLE_HC_SMALL_TABLE_XTR_BIT_SIZE 9
`define CREOLE_HC_MAX_ENCODE_TOT_WIDTH 165
`define CREOLE_HC_MAX_SHORT_PER_XFER 4
`define CREOLE_HC_MAX_SHORT_64K 575
`define CREOLE_HC_MAX_LONG_64K  247
`define CREOLE_HC_MAX_SHORT_16K 543
`define CREOLE_HC_MAX_LONG_16K  245
`define CREOLE_HC_MAX_SHORT_8K  527
`define CREOLE_HC_MAX_LONG_8K   244
`define CREOLE_HC_MAX_SHORT_4K  511
`define CREOLE_HC_MAX_LONG_4K   243
`define CREOLE_HC_MAX_LEN_DF    258
`define CREOLE_HC_MAX_DST_DF    32768
`define CREOLE_HC_STCL_MAX_BITS 2**7
`define CREOLE_HC_ST_MAX_BITS   2**13
`define CREOLE_HC_SYMB_MAX_BITS 2**20
`define CREOLE_HC_SYMB_MAX_BITS_WIDTH $clog2(`CREOLE_HC_SYMB_MAX_BITS)
`define CREOLE_HC_STCL_MAX_BITS_WIDTH $clog2(`CREOLE_HC_STCL_MAX_BITS)
`define CREOLE_HC_ST_MAX_BITS_WIDTH $clog2(`CREOLE_HC_ST_MAX_BITS)
`define CREOLE_HC_STCL_ADDR_WIDTH $clog2(`CREOLE_HC_STCL_MAX_BITS/`CREOLE_HC_HDR_WIDTH)
`define CREOLE_HC_ST_ADDR_WIDTH   $clog2(`CREOLE_HC_ST_MAX_BITS/`CREOLE_HC_HDR_WIDTH)
`define CREOLE_HC_ST_TBL_ENTRIES   `CREOLE_HC_ST_MAX_BITS/`CREOLE_HC_HDR_WIDTH
`define CREOLE_HC_STCL_TBL_ENTRIES `CREOLE_HC_STCL_MAX_BITS/`CREOLE_HC_HDR_WIDTH
`define CREOLE_HC_SYM_ENTRY_CNT_WIDTH 15
`define CREOLE_HC_HLIT_WIDTH  5
`define CREOLE_HC_HDIST_WIDTH 5
`define CREOLE_HC_HCLEN_WIDTH 4
`define CREOLE_HC_LAST_SHORT_PDH 47
`define CREOLE_HC_LAST_LONG_PDH 69
`define CREOLE_HC_BITS_WIDTH 21
`define PRE_HUF_TABLE_NUM_SYM_PER_READ 4
`define MAX_XP_CODE_LENGTH 27
`define HT_FREQ_RD_LATENCY 1
`define MAX_DEFLATE_CODE_LENGTH 15
`define MAX_NUM_SYM_TABLE 704
`define MIN_LITERAL_SYMBOL 257
`define MIN_DISTANCE_SYMBOL 1
`define CREOLE_HC_ST_SYMB_WIDTH 6
`define CREOLE_HC_ST_SYMB_DEPTH 33
`define CREOLE_HC_ST_SYMB_ADDR_WIDTH $clog2(`CREOLE_HC_ST_SYMB_DEPTH)
`define CREOLE_HC_ST_SYMB_FREQ_WIDTH 10
`define CREOLE_HC_MAX_ST_XP_CODE_LENGTH 8
`define CREOLE_HC_MAX_ST_DEFLATE_CODE_LENGTH 7
`define CREOLE_HC_MAX_ST_TABLE_SIZE 33
`define ST_HW_FREQ_RD_LATENCY 2
`define CREOLE_HC_SYM_CODELENGTH $clog2(`MAX_XP_CODE_LENGTH+1)
`define CREOLE_HC_ST_SYM_CODELENGTH $clog2(`CREOLE_HC_MAX_ST_XP_CODE_LENGTH+1)
`define MAX_SHORT_ST_ENTRIES_USED 584
`define MAX_LONG_ST_ENTRIES_USED 249

`define HE_XP_FILL_CNT 16
`define HE_XP_FILL_ENCODE 6'd28
`define HE_XP_ZR_RPT_ENCODE 6'd29
`define HE_XP_PREV_ENCODE 6'd30
`define HE_XP_ROW_0_ENCODE 6'd31
`define HE_XP_ROW_1_ENCODE 6'd32

`define HE_DFLT_LO_ZR_RPT_THRESHOLD 3
`define HE_DFLT_HI_ZR_RPT_THRESHOLD 11
`define HE_DFLT_MX_ZR_RPT_THRESHOLD 138
`define HE_DFLT_NZ_RPT_SYM 16
`define HE_DFLT_LO_NZ_RPT_THRESHOLD 3
`define HE_DFLT_HI_NZ_RPT_THRESHOLD 6
`define HE_DFLT_LO_ZR_RPT_SYM 17
`define HE_DFLT_HI_ZR_RPT_SYM 18
  
`include "cr_huf_compPKG.svp"
`endif 



    

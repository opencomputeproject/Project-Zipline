/*************************************************************************
*
* Copyright © Microsoft Corporation. All rights reserved.
* Copyright © Broadcom Inc. All rights reserved.
* Licensed under the MIT License.
*
*************************************************************************/

`define CR_BIMC_MONITOR_T_DECL   31:0
`define CR_BIMC_MONITOR_T_WIDTH  32
  `define CR_BIMC_MONITOR_T_DEFAULT  (32'h 0)

`define CR_BIMC_MONITOR_T_UNCORRECTABLE_ECC_ERROR_DECL   0:0
`define CR_BIMC_MONITOR_T_UNCORRECTABLE_ECC_ERROR_WIDTH  1
  `define CR_BIMC_MONITOR_T_UNCORRECTABLE_ECC_ERROR_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_T_CORRECTABLE_ECC_ERROR_DECL   0:0
`define CR_BIMC_MONITOR_T_CORRECTABLE_ECC_ERROR_WIDTH  1
  `define CR_BIMC_MONITOR_T_CORRECTABLE_ECC_ERROR_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_T_PARITY_ERROR_DECL   0:0
`define CR_BIMC_MONITOR_T_PARITY_ERROR_WIDTH  1
  `define CR_BIMC_MONITOR_T_PARITY_ERROR_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_T_RESERVE_DECL   0:0
`define CR_BIMC_MONITOR_T_RESERVE_WIDTH  1
  `define CR_BIMC_MONITOR_T_RESERVE_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_T_BIMC_CHAIN_RCV_ERROR_DECL   0:0
`define CR_BIMC_MONITOR_T_BIMC_CHAIN_RCV_ERROR_WIDTH  1
  `define CR_BIMC_MONITOR_T_BIMC_CHAIN_RCV_ERROR_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_T_RCV_INVALID_OPCODE_DECL   0:0
`define CR_BIMC_MONITOR_T_RCV_INVALID_OPCODE_WIDTH  1
  `define CR_BIMC_MONITOR_T_RCV_INVALID_OPCODE_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_T_UNANSWERED_READ_DECL   0:0
`define CR_BIMC_MONITOR_T_UNANSWERED_READ_WIDTH  1
  `define CR_BIMC_MONITOR_T_UNANSWERED_READ_DEFAULT  (1'h 0)

`define CR_FULL_BIMC_MONITOR_T_DECL   31:0
`define CR_FULL_BIMC_MONITOR_T_WIDTH  32
  `define CR_FULL_BIMC_MONITOR_T_UNCORRECTABLE_ECC_ERROR  0
  `define CR_FULL_BIMC_MONITOR_T_CORRECTABLE_ECC_ERROR    1
  `define CR_FULL_BIMC_MONITOR_T_PARITY_ERROR             2
  `define CR_FULL_BIMC_MONITOR_T_RESERVE                  3
  `define CR_FULL_BIMC_MONITOR_T_BIMC_CHAIN_RCV_ERROR     4
  `define CR_FULL_BIMC_MONITOR_T_RCV_INVALID_OPCODE       5
  `define CR_FULL_BIMC_MONITOR_T_UNANSWERED_READ          6
  `define CR_FULL_BIMC_MONITOR_T_RESERVED0                31:7

`define CR_C_BIMC_MONITOR_T_DECL   6:0
`define CR_C_BIMC_MONITOR_T_WIDTH  7
  `define CR_C_BIMC_MONITOR_T_UNCORRECTABLE_ECC_ERROR  0
  `define CR_C_BIMC_MONITOR_T_CORRECTABLE_ECC_ERROR    1
  `define CR_C_BIMC_MONITOR_T_PARITY_ERROR             2
  `define CR_C_BIMC_MONITOR_T_RESERVE                  3
  `define CR_C_BIMC_MONITOR_T_BIMC_CHAIN_RCV_ERROR     4
  `define CR_C_BIMC_MONITOR_T_RCV_INVALID_OPCODE       5
  `define CR_C_BIMC_MONITOR_T_UNANSWERED_READ          6

`define CR_BIMC_MONITOR_MASK_T_DECL   31:0
`define CR_BIMC_MONITOR_MASK_T_WIDTH  32
  `define CR_BIMC_MONITOR_MASK_T_DEFAULT  (32'h 0)

`define CR_BIMC_MONITOR_MASK_T_UNCORRECTABLE_ECC_ERROR_ENABLE_DECL   0:0
`define CR_BIMC_MONITOR_MASK_T_UNCORRECTABLE_ECC_ERROR_ENABLE_WIDTH  1
  `define CR_BIMC_MONITOR_MASK_T_UNCORRECTABLE_ECC_ERROR_ENABLE_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_MASK_T_CORRECTABLE_ECC_ERROR_ENABLE_DECL   0:0
`define CR_BIMC_MONITOR_MASK_T_CORRECTABLE_ECC_ERROR_ENABLE_WIDTH  1
  `define CR_BIMC_MONITOR_MASK_T_CORRECTABLE_ECC_ERROR_ENABLE_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_MASK_T_PARITY_ERROR_ENABLE_DECL   0:0
`define CR_BIMC_MONITOR_MASK_T_PARITY_ERROR_ENABLE_WIDTH  1
  `define CR_BIMC_MONITOR_MASK_T_PARITY_ERROR_ENABLE_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_MASK_T_RESERVE_DECL   0:0
`define CR_BIMC_MONITOR_MASK_T_RESERVE_WIDTH  1
  `define CR_BIMC_MONITOR_MASK_T_RESERVE_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_MASK_T_BIMC_CHAIN_RCV_ERROR_ENABLE_DECL   0:0
`define CR_BIMC_MONITOR_MASK_T_BIMC_CHAIN_RCV_ERROR_ENABLE_WIDTH  1
  `define CR_BIMC_MONITOR_MASK_T_BIMC_CHAIN_RCV_ERROR_ENABLE_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_MASK_T_RCV_INVALID_OPCODE_DECL   0:0
`define CR_BIMC_MONITOR_MASK_T_RCV_INVALID_OPCODE_WIDTH  1
  `define CR_BIMC_MONITOR_MASK_T_RCV_INVALID_OPCODE_DEFAULT  (1'h 0)

`define CR_BIMC_MONITOR_MASK_T_UNANSWERED_READ_DECL   0:0
`define CR_BIMC_MONITOR_MASK_T_UNANSWERED_READ_WIDTH  1
  `define CR_BIMC_MONITOR_MASK_T_UNANSWERED_READ_DEFAULT  (1'h 0)

`define CR_FULL_BIMC_MONITOR_MASK_T_DECL   31:0
`define CR_FULL_BIMC_MONITOR_MASK_T_WIDTH  32
  `define CR_FULL_BIMC_MONITOR_MASK_T_UNCORRECTABLE_ECC_ERROR_ENABLE  0
  `define CR_FULL_BIMC_MONITOR_MASK_T_CORRECTABLE_ECC_ERROR_ENABLE    1
  `define CR_FULL_BIMC_MONITOR_MASK_T_PARITY_ERROR_ENABLE             2
  `define CR_FULL_BIMC_MONITOR_MASK_T_RESERVE                         3
  `define CR_FULL_BIMC_MONITOR_MASK_T_BIMC_CHAIN_RCV_ERROR_ENABLE     4
  `define CR_FULL_BIMC_MONITOR_MASK_T_RCV_INVALID_OPCODE              5
  `define CR_FULL_BIMC_MONITOR_MASK_T_UNANSWERED_READ                 6
  `define CR_FULL_BIMC_MONITOR_MASK_T_RESERVED0                       31:7

`define CR_C_BIMC_MONITOR_MASK_T_DECL   6:0
`define CR_C_BIMC_MONITOR_MASK_T_WIDTH  7
  `define CR_C_BIMC_MONITOR_MASK_T_UNCORRECTABLE_ECC_ERROR_ENABLE  0
  `define CR_C_BIMC_MONITOR_MASK_T_CORRECTABLE_ECC_ERROR_ENABLE    1
  `define CR_C_BIMC_MONITOR_MASK_T_PARITY_ERROR_ENABLE             2
  `define CR_C_BIMC_MONITOR_MASK_T_RESERVE                         3
  `define CR_C_BIMC_MONITOR_MASK_T_BIMC_CHAIN_RCV_ERROR_ENABLE     4
  `define CR_C_BIMC_MONITOR_MASK_T_RCV_INVALID_OPCODE              5
  `define CR_C_BIMC_MONITOR_MASK_T_UNANSWERED_READ                 6

`define CR_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_DECL   31:0
`define CR_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_WIDTH  32
  `define CR_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_DEFAULT  (32'h 0)

`define CR_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_UNCORRECTABLE_ECC_DECL   31:0
`define CR_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_UNCORRECTABLE_ECC_WIDTH  32
  `define CR_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_UNCORRECTABLE_ECC_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_DECL   31:0
`define CR_FULL_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_WIDTH  32
  `define CR_FULL_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_UNCORRECTABLE_ECC  31:00

`define CR_C_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_DECL   31:0
`define CR_C_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_WIDTH  32
  `define CR_C_BIMC_ECC_UNCORRECTABLE_ERROR_CNT_T_UNCORRECTABLE_ECC  31:00

`define CR_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_DECL   31:0
`define CR_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_WIDTH  32
  `define CR_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_DEFAULT  (32'h 0)

`define CR_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_CORRECTABLE_ECC_DECL   31:0
`define CR_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_CORRECTABLE_ECC_WIDTH  32
  `define CR_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_CORRECTABLE_ECC_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_DECL   31:0
`define CR_FULL_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_WIDTH  32
  `define CR_FULL_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_CORRECTABLE_ECC  31:00

`define CR_C_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_DECL   31:0
`define CR_C_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_WIDTH  32
  `define CR_C_BIMC_ECC_CORRECTABLE_ERROR_CNT_T_CORRECTABLE_ECC  31:00

`define CR_BIMC_PARITY_ERROR_CNT_T_DECL   31:0
`define CR_BIMC_PARITY_ERROR_CNT_T_WIDTH  32
  `define CR_BIMC_PARITY_ERROR_CNT_T_DEFAULT  (32'h 0)

`define CR_BIMC_PARITY_ERROR_CNT_T_PARITY_ERRORS_DECL   31:0
`define CR_BIMC_PARITY_ERROR_CNT_T_PARITY_ERRORS_WIDTH  32
  `define CR_BIMC_PARITY_ERROR_CNT_T_PARITY_ERRORS_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_PARITY_ERROR_CNT_T_DECL   31:0
`define CR_FULL_BIMC_PARITY_ERROR_CNT_T_WIDTH  32
  `define CR_FULL_BIMC_PARITY_ERROR_CNT_T_PARITY_ERRORS  31:00

`define CR_C_BIMC_PARITY_ERROR_CNT_T_DECL   31:0
`define CR_C_BIMC_PARITY_ERROR_CNT_T_WIDTH  32
  `define CR_C_BIMC_PARITY_ERROR_CNT_T_PARITY_ERRORS  31:00

`define CR_BIMC_GLOBAL_CONFIG_T_DECL   31:0
`define CR_BIMC_GLOBAL_CONFIG_T_WIDTH  32
  `define CR_BIMC_GLOBAL_CONFIG_T_DEFAULT  (32'h 1)

`define CR_BIMC_GLOBAL_CONFIG_T_SOFT_RESET_DECL   0:0
`define CR_BIMC_GLOBAL_CONFIG_T_SOFT_RESET_WIDTH  1
  `define CR_BIMC_GLOBAL_CONFIG_T_SOFT_RESET_DEFAULT  (1'h 1)

`define CR_BIMC_GLOBAL_CONFIG_T_RESERVE_DECL   0:0
`define CR_BIMC_GLOBAL_CONFIG_T_RESERVE_WIDTH  1
  `define CR_BIMC_GLOBAL_CONFIG_T_RESERVE_DEFAULT  (1'h 0)

`define CR_BIMC_GLOBAL_CONFIG_T_BIMC_MEM_INIT_DONE_DECL   0:0
`define CR_BIMC_GLOBAL_CONFIG_T_BIMC_MEM_INIT_DONE_WIDTH  1
  `define CR_BIMC_GLOBAL_CONFIG_T_BIMC_MEM_INIT_DONE_DEFAULT  (1'h 0)

`define CR_BIMC_GLOBAL_CONFIG_T_MEM_WR_INIT_DECL   0:0
`define CR_BIMC_GLOBAL_CONFIG_T_MEM_WR_INIT_WIDTH  1
  `define CR_BIMC_GLOBAL_CONFIG_T_MEM_WR_INIT_DEFAULT  (1'h 0)

`define CR_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_ERROR_DECL   0:0
`define CR_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_ERROR_WIDTH  1
  `define CR_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_ERROR_DEFAULT  (1'h 0)

`define CR_BIMC_GLOBAL_CONFIG_T_DEBUG_WRITE_EN_DECL   0:0
`define CR_BIMC_GLOBAL_CONFIG_T_DEBUG_WRITE_EN_WIDTH  1
  `define CR_BIMC_GLOBAL_CONFIG_T_DEBUG_WRITE_EN_DEFAULT  (1'h 0)

`define CR_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_TIMER_DECL   25:0
`define CR_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_TIMER_WIDTH  26
  `define CR_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_TIMER_DEFAULT  (26'h 0)

`define CR_FULL_BIMC_GLOBAL_CONFIG_T_DECL   31:0
`define CR_FULL_BIMC_GLOBAL_CONFIG_T_WIDTH  32
  `define CR_FULL_BIMC_GLOBAL_CONFIG_T_SOFT_RESET          00
  `define CR_FULL_BIMC_GLOBAL_CONFIG_T_RESERVE             01
  `define CR_FULL_BIMC_GLOBAL_CONFIG_T_BIMC_MEM_INIT_DONE  02
  `define CR_FULL_BIMC_GLOBAL_CONFIG_T_MEM_WR_INIT         03
  `define CR_FULL_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_ERROR  04
  `define CR_FULL_BIMC_GLOBAL_CONFIG_T_DEBUG_WRITE_EN      05
  `define CR_FULL_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_TIMER  31:06

`define CR_C_BIMC_GLOBAL_CONFIG_T_DECL   31:0
`define CR_C_BIMC_GLOBAL_CONFIG_T_WIDTH  32
  `define CR_C_BIMC_GLOBAL_CONFIG_T_SOFT_RESET          00
  `define CR_C_BIMC_GLOBAL_CONFIG_T_RESERVE             01
  `define CR_C_BIMC_GLOBAL_CONFIG_T_BIMC_MEM_INIT_DONE  02
  `define CR_C_BIMC_GLOBAL_CONFIG_T_MEM_WR_INIT         03
  `define CR_C_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_ERROR  04
  `define CR_C_BIMC_GLOBAL_CONFIG_T_DEBUG_WRITE_EN      05
  `define CR_C_BIMC_GLOBAL_CONFIG_T_POLL_ECC_PAR_TIMER  31:06

`define CR_BIMC_MEMID_T_DECL   31:0
`define CR_BIMC_MEMID_T_WIDTH  32
  `define CR_BIMC_MEMID_T_DEFAULT  (32'h 0)

`define CR_BIMC_MEMID_T_MAX_MEMID_DECL   11:0
`define CR_BIMC_MEMID_T_MAX_MEMID_WIDTH  12
  `define CR_BIMC_MEMID_T_MAX_MEMID_DEFAULT  (12'h 0)

`define CR_FULL_BIMC_MEMID_T_DECL   31:0
`define CR_FULL_BIMC_MEMID_T_WIDTH  32
  `define CR_FULL_BIMC_MEMID_T_MAX_MEMID  11:00
  `define CR_FULL_BIMC_MEMID_T_RESERVED0  31:12

`define CR_C_BIMC_MEMID_T_DECL   11:0
`define CR_C_BIMC_MEMID_T_WIDTH  12
  `define CR_C_BIMC_MEMID_T_MAX_MEMID  11:00

`define CR_BIMC_ECCPAR_DEBUG_T_DECL   31:0
`define CR_BIMC_ECCPAR_DEBUG_T_WIDTH  32
  `define CR_BIMC_ECCPAR_DEBUG_T_DEFAULT  (32'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_MEMADDR_DECL   11:0
`define CR_BIMC_ECCPAR_DEBUG_T_MEMADDR_WIDTH  12
  `define CR_BIMC_ECCPAR_DEBUG_T_MEMADDR_DEFAULT  (12'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_MEMTYPE_DECL   3:0
`define CR_BIMC_ECCPAR_DEBUG_T_MEMTYPE_WIDTH  4
  `define CR_BIMC_ECCPAR_DEBUG_T_MEMTYPE_DEFAULT  (4'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_ECCPAR_CORRUPT_DECL   1:0
`define CR_BIMC_ECCPAR_DEBUG_T_ECCPAR_CORRUPT_WIDTH  2
  `define CR_BIMC_ECCPAR_DEBUG_T_ECCPAR_CORRUPT_DEFAULT  (2'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_RESERVE_DECL   1:0
`define CR_BIMC_ECCPAR_DEBUG_T_RESERVE_WIDTH  2
  `define CR_BIMC_ECCPAR_DEBUG_T_RESERVE_DEFAULT  (2'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_ECCPAR_DISABLE_DECL   1:0
`define CR_BIMC_ECCPAR_DEBUG_T_ECCPAR_DISABLE_WIDTH  2
  `define CR_BIMC_ECCPAR_DEBUG_T_ECCPAR_DISABLE_DEFAULT  (2'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_SEND_DECL   0:0
`define CR_BIMC_ECCPAR_DEBUG_T_SEND_WIDTH  1
  `define CR_BIMC_ECCPAR_DEBUG_T_SEND_DEFAULT  (1'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_SENT_DECL   0:0
`define CR_BIMC_ECCPAR_DEBUG_T_SENT_WIDTH  1
  `define CR_BIMC_ECCPAR_DEBUG_T_SENT_DEFAULT  (1'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_JABBER_OFF_DECL   3:0
`define CR_BIMC_ECCPAR_DEBUG_T_JABBER_OFF_WIDTH  4
  `define CR_BIMC_ECCPAR_DEBUG_T_JABBER_OFF_DEFAULT  (4'h 0)

`define CR_BIMC_ECCPAR_DEBUG_T_ACK_DECL   0:0
`define CR_BIMC_ECCPAR_DEBUG_T_ACK_WIDTH  1
  `define CR_BIMC_ECCPAR_DEBUG_T_ACK_DEFAULT  (1'h 0)

`define CR_FULL_BIMC_ECCPAR_DEBUG_T_DECL   31:0
`define CR_FULL_BIMC_ECCPAR_DEBUG_T_WIDTH  32
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_MEMADDR         11:00
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_MEMTYPE         15:12
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_ECCPAR_CORRUPT  17:16
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_RESERVE         19:18
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_ECCPAR_DISABLE  21:20
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_SEND            22
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_SENT            23
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_JABBER_OFF      27:24
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_ACK             28
  `define CR_FULL_BIMC_ECCPAR_DEBUG_T_RESERVED0       31:29

`define CR_C_BIMC_ECCPAR_DEBUG_T_DECL   28:0
`define CR_C_BIMC_ECCPAR_DEBUG_T_WIDTH  29
  `define CR_C_BIMC_ECCPAR_DEBUG_T_MEMADDR         11:00
  `define CR_C_BIMC_ECCPAR_DEBUG_T_MEMTYPE         15:12
  `define CR_C_BIMC_ECCPAR_DEBUG_T_ECCPAR_CORRUPT  17:16
  `define CR_C_BIMC_ECCPAR_DEBUG_T_RESERVE         19:18
  `define CR_C_BIMC_ECCPAR_DEBUG_T_ECCPAR_DISABLE  21:20
  `define CR_C_BIMC_ECCPAR_DEBUG_T_SEND            22
  `define CR_C_BIMC_ECCPAR_DEBUG_T_SENT            23
  `define CR_C_BIMC_ECCPAR_DEBUG_T_JABBER_OFF      27:24
  `define CR_C_BIMC_ECCPAR_DEBUG_T_ACK             28

`define CR_BIMC_CMD2_T_DECL   31:0
`define CR_BIMC_CMD2_T_WIDTH  32
  `define CR_BIMC_CMD2_T_DEFAULT  (32'h 0)

`define CR_BIMC_CMD2_T_OPCODE_DECL   7:0
`define CR_BIMC_CMD2_T_OPCODE_WIDTH  8
  `define CR_BIMC_CMD2_T_OPCODE_DEFAULT  (8'h 0)

`define CR_BIMC_CMD2_T_SEND_DECL   0:0
`define CR_BIMC_CMD2_T_SEND_WIDTH  1
  `define CR_BIMC_CMD2_T_SEND_DEFAULT  (1'h 0)

`define CR_BIMC_CMD2_T_SENT_DECL   0:0
`define CR_BIMC_CMD2_T_SENT_WIDTH  1
  `define CR_BIMC_CMD2_T_SENT_DEFAULT  (1'h 0)

`define CR_BIMC_CMD2_T_ACK_DECL   0:0
`define CR_BIMC_CMD2_T_ACK_WIDTH  1
  `define CR_BIMC_CMD2_T_ACK_DEFAULT  (1'h 0)

`define CR_FULL_BIMC_CMD2_T_DECL   31:0
`define CR_FULL_BIMC_CMD2_T_WIDTH  32
  `define CR_FULL_BIMC_CMD2_T_OPCODE     07:00
  `define CR_FULL_BIMC_CMD2_T_SEND       08
  `define CR_FULL_BIMC_CMD2_T_SENT       09
  `define CR_FULL_BIMC_CMD2_T_ACK        10
  `define CR_FULL_BIMC_CMD2_T_RESERVED0  31:11

`define CR_C_BIMC_CMD2_T_DECL   10:0
`define CR_C_BIMC_CMD2_T_WIDTH  11
  `define CR_C_BIMC_CMD2_T_OPCODE  07:00
  `define CR_C_BIMC_CMD2_T_SEND    08
  `define CR_C_BIMC_CMD2_T_SENT    09
  `define CR_C_BIMC_CMD2_T_ACK     10

`define CR_BIMC_CMD1_T_DECL   31:0
`define CR_BIMC_CMD1_T_WIDTH  32
  `define CR_BIMC_CMD1_T_DEFAULT  (32'h 0)

`define CR_BIMC_CMD1_T_ADDR_DECL   15:0
`define CR_BIMC_CMD1_T_ADDR_WIDTH  16
  `define CR_BIMC_CMD1_T_ADDR_DEFAULT  (16'h 0)

`define CR_BIMC_CMD1_T_MEM_DECL   11:0
`define CR_BIMC_CMD1_T_MEM_WIDTH  12
  `define CR_BIMC_CMD1_T_MEM_DEFAULT  (12'h 0)

`define CR_BIMC_CMD1_T_MEMTYPE_DECL   3:0
`define CR_BIMC_CMD1_T_MEMTYPE_WIDTH  4
  `define CR_BIMC_CMD1_T_MEMTYPE_DEFAULT  (4'h 0)

`define CR_FULL_BIMC_CMD1_T_DECL   31:0
`define CR_FULL_BIMC_CMD1_T_WIDTH  32
  `define CR_FULL_BIMC_CMD1_T_ADDR     15:00
  `define CR_FULL_BIMC_CMD1_T_MEM      27:16
  `define CR_FULL_BIMC_CMD1_T_MEMTYPE  31:28

`define CR_C_BIMC_CMD1_T_DECL   31:0
`define CR_C_BIMC_CMD1_T_WIDTH  32
  `define CR_C_BIMC_CMD1_T_ADDR     15:00
  `define CR_C_BIMC_CMD1_T_MEM      27:16
  `define CR_C_BIMC_CMD1_T_MEMTYPE  31:28

`define CR_BIMC_CMD0_T_DECL   31:0
`define CR_BIMC_CMD0_T_WIDTH  32
  `define CR_BIMC_CMD0_T_DEFAULT  (32'h 0)

`define CR_BIMC_CMD0_T_DATA_DECL   31:0
`define CR_BIMC_CMD0_T_DATA_WIDTH  32
  `define CR_BIMC_CMD0_T_DATA_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_CMD0_T_DECL   31:0
`define CR_FULL_BIMC_CMD0_T_WIDTH  32
  `define CR_FULL_BIMC_CMD0_T_DATA  31:00

`define CR_C_BIMC_CMD0_T_DECL   31:0
`define CR_C_BIMC_CMD0_T_WIDTH  32
  `define CR_C_BIMC_CMD0_T_DATA  31:00

`define CR_BIMC_RXCMD2_T_DECL   31:0
`define CR_BIMC_RXCMD2_T_WIDTH  32
  `define CR_BIMC_RXCMD2_T_DEFAULT  (32'h 0)

`define CR_BIMC_RXCMD2_T_OPCODE_DECL   7:0
`define CR_BIMC_RXCMD2_T_OPCODE_WIDTH  8
  `define CR_BIMC_RXCMD2_T_OPCODE_DEFAULT  (8'h 0)

`define CR_BIMC_RXCMD2_T_RXFLAG_DECL   0:0
`define CR_BIMC_RXCMD2_T_RXFLAG_WIDTH  1
  `define CR_BIMC_RXCMD2_T_RXFLAG_DEFAULT  (1'h 0)

`define CR_BIMC_RXCMD2_T_ACK_DECL   0:0
`define CR_BIMC_RXCMD2_T_ACK_WIDTH  1

`define CR_FULL_BIMC_RXCMD2_T_DECL   31:0
`define CR_FULL_BIMC_RXCMD2_T_WIDTH  32
  `define CR_FULL_BIMC_RXCMD2_T_OPCODE     7:0
  `define CR_FULL_BIMC_RXCMD2_T_RXFLAG     8
  `define CR_FULL_BIMC_RXCMD2_T_ACK        9
  `define CR_FULL_BIMC_RXCMD2_T_RESERVED0  31:10

`define CR_C_BIMC_RXCMD2_T_DECL   9:0
`define CR_C_BIMC_RXCMD2_T_WIDTH  10
  `define CR_C_BIMC_RXCMD2_T_OPCODE  7:0
  `define CR_C_BIMC_RXCMD2_T_RXFLAG  8
  `define CR_C_BIMC_RXCMD2_T_ACK     9

`define CR_BIMC_RXCMD1_T_DECL   31:0
`define CR_BIMC_RXCMD1_T_WIDTH  32
  `define CR_BIMC_RXCMD1_T_DEFAULT  (32'h 0)

`define CR_BIMC_RXCMD1_T_ADDR_DECL   15:0
`define CR_BIMC_RXCMD1_T_ADDR_WIDTH  16
  `define CR_BIMC_RXCMD1_T_ADDR_DEFAULT  (16'h 0)

`define CR_BIMC_RXCMD1_T_MEM_DECL   11:0
`define CR_BIMC_RXCMD1_T_MEM_WIDTH  12
  `define CR_BIMC_RXCMD1_T_MEM_DEFAULT  (12'h 0)

`define CR_BIMC_RXCMD1_T_MEMTYPE_DECL   3:0
`define CR_BIMC_RXCMD1_T_MEMTYPE_WIDTH  4
  `define CR_BIMC_RXCMD1_T_MEMTYPE_DEFAULT  (4'h 0)

`define CR_FULL_BIMC_RXCMD1_T_DECL   31:0
`define CR_FULL_BIMC_RXCMD1_T_WIDTH  32
  `define CR_FULL_BIMC_RXCMD1_T_ADDR     15:00
  `define CR_FULL_BIMC_RXCMD1_T_MEM      27:16
  `define CR_FULL_BIMC_RXCMD1_T_MEMTYPE  31:28

`define CR_C_BIMC_RXCMD1_T_DECL   31:0
`define CR_C_BIMC_RXCMD1_T_WIDTH  32
  `define CR_C_BIMC_RXCMD1_T_ADDR     15:00
  `define CR_C_BIMC_RXCMD1_T_MEM      27:16
  `define CR_C_BIMC_RXCMD1_T_MEMTYPE  31:28

`define CR_BIMC_RXCMD0_T_DECL   31:0
`define CR_BIMC_RXCMD0_T_WIDTH  32
  `define CR_BIMC_RXCMD0_T_DEFAULT  (32'h 0)

`define CR_BIMC_RXCMD0_T_DATA_DECL   31:0
`define CR_BIMC_RXCMD0_T_DATA_WIDTH  32
  `define CR_BIMC_RXCMD0_T_DATA_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_RXCMD0_T_DECL   31:0
`define CR_FULL_BIMC_RXCMD0_T_WIDTH  32
  `define CR_FULL_BIMC_RXCMD0_T_DATA  31:00

`define CR_C_BIMC_RXCMD0_T_DECL   31:0
`define CR_C_BIMC_RXCMD0_T_WIDTH  32
  `define CR_C_BIMC_RXCMD0_T_DATA  31:00

`define CR_BIMC_RXRSP2_T_DECL   31:0
`define CR_BIMC_RXRSP2_T_WIDTH  32
  `define CR_BIMC_RXRSP2_T_DEFAULT  (32'h 0)

`define CR_BIMC_RXRSP2_T_DATA_DECL   7:0
`define CR_BIMC_RXRSP2_T_DATA_WIDTH  8
  `define CR_BIMC_RXRSP2_T_DATA_DEFAULT  (8'h 0)

`define CR_BIMC_RXRSP2_T_RXFLAG_DECL   0:0
`define CR_BIMC_RXRSP2_T_RXFLAG_WIDTH  1
  `define CR_BIMC_RXRSP2_T_RXFLAG_DEFAULT  (1'h 0)

`define CR_BIMC_RXRSP2_T_ACK_DECL   0:0
`define CR_BIMC_RXRSP2_T_ACK_WIDTH  1

`define CR_FULL_BIMC_RXRSP2_T_DECL   31:0
`define CR_FULL_BIMC_RXRSP2_T_WIDTH  32
  `define CR_FULL_BIMC_RXRSP2_T_DATA       7:0
  `define CR_FULL_BIMC_RXRSP2_T_RXFLAG     8
  `define CR_FULL_BIMC_RXRSP2_T_ACK        9
  `define CR_FULL_BIMC_RXRSP2_T_RESERVED0  31:10

`define CR_C_BIMC_RXRSP2_T_DECL   9:0
`define CR_C_BIMC_RXRSP2_T_WIDTH  10
  `define CR_C_BIMC_RXRSP2_T_DATA    7:0
  `define CR_C_BIMC_RXRSP2_T_RXFLAG  8
  `define CR_C_BIMC_RXRSP2_T_ACK     9

`define CR_BIMC_RXRSP1_T_DECL   31:0
`define CR_BIMC_RXRSP1_T_WIDTH  32
  `define CR_BIMC_RXRSP1_T_DEFAULT  (32'h 0)

`define CR_BIMC_RXRSP1_T_DATA_DECL   31:0
`define CR_BIMC_RXRSP1_T_DATA_WIDTH  32
  `define CR_BIMC_RXRSP1_T_DATA_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_RXRSP1_T_DECL   31:0
`define CR_FULL_BIMC_RXRSP1_T_WIDTH  32
  `define CR_FULL_BIMC_RXRSP1_T_DATA  31:00

`define CR_C_BIMC_RXRSP1_T_DECL   31:0
`define CR_C_BIMC_RXRSP1_T_WIDTH  32
  `define CR_C_BIMC_RXRSP1_T_DATA  31:00

`define CR_BIMC_RXRSP0_T_DECL   31:0
`define CR_BIMC_RXRSP0_T_WIDTH  32
  `define CR_BIMC_RXRSP0_T_DEFAULT  (32'h 0)

`define CR_BIMC_RXRSP0_T_DATA_DECL   31:0
`define CR_BIMC_RXRSP0_T_DATA_WIDTH  32
  `define CR_BIMC_RXRSP0_T_DATA_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_RXRSP0_T_DECL   31:0
`define CR_FULL_BIMC_RXRSP0_T_WIDTH  32
  `define CR_FULL_BIMC_RXRSP0_T_DATA  31:00

`define CR_C_BIMC_RXRSP0_T_DECL   31:0
`define CR_C_BIMC_RXRSP0_T_WIDTH  32
  `define CR_C_BIMC_RXRSP0_T_DATA  31:00

`define CR_BIMC_POLLRSP2_T_DECL   31:0
`define CR_BIMC_POLLRSP2_T_WIDTH  32
  `define CR_BIMC_POLLRSP2_T_DEFAULT  (32'h 0)

`define CR_BIMC_POLLRSP2_T_DATA_DECL   7:0
`define CR_BIMC_POLLRSP2_T_DATA_WIDTH  8
  `define CR_BIMC_POLLRSP2_T_DATA_DEFAULT  (8'h 0)

`define CR_BIMC_POLLRSP2_T_RXFLAG_DECL   0:0
`define CR_BIMC_POLLRSP2_T_RXFLAG_WIDTH  1
  `define CR_BIMC_POLLRSP2_T_RXFLAG_DEFAULT  (1'h 0)

`define CR_BIMC_POLLRSP2_T_ACK_DECL   0:0
`define CR_BIMC_POLLRSP2_T_ACK_WIDTH  1

`define CR_FULL_BIMC_POLLRSP2_T_DECL   31:0
`define CR_FULL_BIMC_POLLRSP2_T_WIDTH  32
  `define CR_FULL_BIMC_POLLRSP2_T_DATA       7:0
  `define CR_FULL_BIMC_POLLRSP2_T_RXFLAG     8
  `define CR_FULL_BIMC_POLLRSP2_T_ACK        9
  `define CR_FULL_BIMC_POLLRSP2_T_RESERVED0  31:10

`define CR_C_BIMC_POLLRSP2_T_DECL   9:0
`define CR_C_BIMC_POLLRSP2_T_WIDTH  10
  `define CR_C_BIMC_POLLRSP2_T_DATA    7:0
  `define CR_C_BIMC_POLLRSP2_T_RXFLAG  8
  `define CR_C_BIMC_POLLRSP2_T_ACK     9

`define CR_BIMC_POLLRSP1_T_DECL   31:0
`define CR_BIMC_POLLRSP1_T_WIDTH  32
  `define CR_BIMC_POLLRSP1_T_DEFAULT  (32'h 0)

`define CR_BIMC_POLLRSP1_T_DATA_DECL   31:0
`define CR_BIMC_POLLRSP1_T_DATA_WIDTH  32
  `define CR_BIMC_POLLRSP1_T_DATA_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_POLLRSP1_T_DECL   31:0
`define CR_FULL_BIMC_POLLRSP1_T_WIDTH  32
  `define CR_FULL_BIMC_POLLRSP1_T_DATA  31:00

`define CR_C_BIMC_POLLRSP1_T_DECL   31:0
`define CR_C_BIMC_POLLRSP1_T_WIDTH  32
  `define CR_C_BIMC_POLLRSP1_T_DATA  31:00

`define CR_BIMC_POLLRSP0_T_DECL   31:0
`define CR_BIMC_POLLRSP0_T_WIDTH  32
  `define CR_BIMC_POLLRSP0_T_DEFAULT  (32'h 0)

`define CR_BIMC_POLLRSP0_T_DATA_DECL   31:0
`define CR_BIMC_POLLRSP0_T_DATA_WIDTH  32
  `define CR_BIMC_POLLRSP0_T_DATA_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_POLLRSP0_T_DECL   31:0
`define CR_FULL_BIMC_POLLRSP0_T_WIDTH  32
  `define CR_FULL_BIMC_POLLRSP0_T_DATA  31:00

`define CR_C_BIMC_POLLRSP0_T_DECL   31:0
`define CR_C_BIMC_POLLRSP0_T_WIDTH  32
  `define CR_C_BIMC_POLLRSP0_T_DATA  31:00

`define CR_BIMC_DBGCMD2_T_DECL   31:0
`define CR_BIMC_DBGCMD2_T_WIDTH  32
  `define CR_BIMC_DBGCMD2_T_DEFAULT  (32'h 0)

`define CR_BIMC_DBGCMD2_T_OPCODE_DECL   7:0
`define CR_BIMC_DBGCMD2_T_OPCODE_WIDTH  8
  `define CR_BIMC_DBGCMD2_T_OPCODE_DEFAULT  (8'h 0)

`define CR_BIMC_DBGCMD2_T_RXFLAG_DECL   0:0
`define CR_BIMC_DBGCMD2_T_RXFLAG_WIDTH  1
  `define CR_BIMC_DBGCMD2_T_RXFLAG_DEFAULT  (1'h 0)

`define CR_BIMC_DBGCMD2_T_ACK_DECL   0:0
`define CR_BIMC_DBGCMD2_T_ACK_WIDTH  1

`define CR_FULL_BIMC_DBGCMD2_T_DECL   31:0
`define CR_FULL_BIMC_DBGCMD2_T_WIDTH  32
  `define CR_FULL_BIMC_DBGCMD2_T_OPCODE     7:0
  `define CR_FULL_BIMC_DBGCMD2_T_RXFLAG     8
  `define CR_FULL_BIMC_DBGCMD2_T_ACK        9
  `define CR_FULL_BIMC_DBGCMD2_T_RESERVED0  31:10

`define CR_C_BIMC_DBGCMD2_T_DECL   9:0
`define CR_C_BIMC_DBGCMD2_T_WIDTH  10
  `define CR_C_BIMC_DBGCMD2_T_OPCODE  7:0
  `define CR_C_BIMC_DBGCMD2_T_RXFLAG  8
  `define CR_C_BIMC_DBGCMD2_T_ACK     9

`define CR_BIMC_DBGCMD1_T_DECL   31:0
`define CR_BIMC_DBGCMD1_T_WIDTH  32
  `define CR_BIMC_DBGCMD1_T_DEFAULT  (32'h 0)

`define CR_BIMC_DBGCMD1_T_ADDR_DECL   15:0
`define CR_BIMC_DBGCMD1_T_ADDR_WIDTH  16
  `define CR_BIMC_DBGCMD1_T_ADDR_DEFAULT  (16'h 0)

`define CR_BIMC_DBGCMD1_T_MEM_DECL   11:0
`define CR_BIMC_DBGCMD1_T_MEM_WIDTH  12
  `define CR_BIMC_DBGCMD1_T_MEM_DEFAULT  (12'h 0)

`define CR_BIMC_DBGCMD1_T_MEMTYPE_DECL   3:0
`define CR_BIMC_DBGCMD1_T_MEMTYPE_WIDTH  4
  `define CR_BIMC_DBGCMD1_T_MEMTYPE_DEFAULT  (4'h 0)

`define CR_FULL_BIMC_DBGCMD1_T_DECL   31:0
`define CR_FULL_BIMC_DBGCMD1_T_WIDTH  32
  `define CR_FULL_BIMC_DBGCMD1_T_ADDR     15:00
  `define CR_FULL_BIMC_DBGCMD1_T_MEM      27:16
  `define CR_FULL_BIMC_DBGCMD1_T_MEMTYPE  31:28

`define CR_C_BIMC_DBGCMD1_T_DECL   31:0
`define CR_C_BIMC_DBGCMD1_T_WIDTH  32
  `define CR_C_BIMC_DBGCMD1_T_ADDR     15:00
  `define CR_C_BIMC_DBGCMD1_T_MEM      27:16
  `define CR_C_BIMC_DBGCMD1_T_MEMTYPE  31:28

`define CR_BIMC_DBGCMD0_T_DECL   31:0
`define CR_BIMC_DBGCMD0_T_WIDTH  32
  `define CR_BIMC_DBGCMD0_T_DEFAULT  (32'h 0)

`define CR_BIMC_DBGCMD0_T_DATA_DECL   31:0
`define CR_BIMC_DBGCMD0_T_DATA_WIDTH  32
  `define CR_BIMC_DBGCMD0_T_DATA_DEFAULT  (32'h 0)

`define CR_FULL_BIMC_DBGCMD0_T_DECL   31:0
`define CR_FULL_BIMC_DBGCMD0_T_WIDTH  32
  `define CR_FULL_BIMC_DBGCMD0_T_DATA  31:00

`define CR_C_BIMC_DBGCMD0_T_DECL   31:0
`define CR_C_BIMC_DBGCMD0_T_WIDTH  32
  `define CR_C_BIMC_DBGCMD0_T_DATA  31:00

  `define CR_BIMC_MONITOR                      ('h 0)
  `define CR_BIMC_MONITOR_MASK                 ('h 4)
  `define CR_BIMC_ECC_UNCORRECTABLE_ERROR_CNT  ('h 8)
  `define CR_BIMC_ECC_CORRECTABLE_ERROR_CNT    ('h c)
  `define CR_BIMC_PARITY_ERROR_CNT             ('h 10)
  `define CR_BIMC_GLOBAL_CONFIG                ('h 14)
  `define CR_BIMC_MEMID                        ('h 18)
  `define CR_BIMC_ECCPAR_DEBUG                 ('h 1c)
  `define CR_BIMC_CMD2                         ('h 20)
  `define CR_BIMC_CMD1                         ('h 24)
  `define CR_BIMC_CMD0                         ('h 28)
  `define CR_BIMC_RXCMD2                       ('h 2c)
  `define CR_BIMC_RXCMD1                       ('h 30)
  `define CR_BIMC_RXCMD0                       ('h 34)
  `define CR_BIMC_RXRSP2                       ('h 38)
  `define CR_BIMC_RXRSP1                       ('h 3c)
  `define CR_BIMC_RXRSP0                       ('h 40)
  `define CR_BIMC_POLLRSP2                     ('h 44)
  `define CR_BIMC_POLLRSP1                     ('h 48)
  `define CR_BIMC_POLLRSP0                     ('h 4c)
  `define CR_BIMC_DBGCMD2                      ('h 50)
  `define CR_BIMC_DBGCMD1                      ('h 54)
  `define CR_BIMC_DBGCMD0                      ('h 58)
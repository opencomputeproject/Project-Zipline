/*************************************************************************
*
* Copyright � Microsoft Corporation. All rights reserved.
* Copyright � Broadcom Inc. All rights reserved.
* Licensed under the MIT License.
*
*************************************************************************/
`define AXI_RS_FULL   0
`define AXI_RS_FWD    1
`define AXI_RS_REV    2
`define AXI_RS_BYPASS 3
/*************************************************************************
*
* Copyright � Microsoft Corporation. All rights reserved.
* Copyright � Broadcom Inc. All rights reserved.
* Licensed under the MIT License.
*
*************************************************************************/








`ifndef __CR_LZ77_COMP_PKG_INCLUDES_VH
`define __CR_LZ77_COMP_PKG_INCLUDES_VH

`include "cr_lz77_comp_regfilePKG.svp"
`include "cr_lz77_comp_regsPKG.svp"
`include "cr_lz77_compPKG.svp"

`endif


/*************************************************************************
*
* Copyright � Microsoft Corporation. All rights reserved.
* Copyright � Broadcom Inc. All rights reserved.
* Licensed under the MIT License.
*
*************************************************************************/








import cr_lz77_compPKG::*;
import cr_lz77_comp_regfilePKG::*;


